module T01(
  input A,B,C,
  output Y);



endmodule
