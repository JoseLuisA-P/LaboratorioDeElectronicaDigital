///////////////////////////////////////////////////////////////////////////////
//Jose Luis Alvarez Pineda
//19392
//Electronica digital
// Muxes para el laboratorio 5
///////////////////////////////////////////////////////////////////////////////
module testbench();

  reg A1,B1,C1;
  wire y;

  //MUX 2:1 de la tabla01
  MUX2T1 sel21(y, A1, B1, C1);

endmodule
