///////////////////////////////////////////////////////////////////////////////
//Jose Luis Alvarez Pineda
//19392
//Electronica digital
// Muxes para el laboratorio 5
///////////////////////////////////////////////////////////////////////////////

//MUX 2:1 de uso general para la practica
module Mux2(
  input wire A,B,S,
  output wire Y);

end module
